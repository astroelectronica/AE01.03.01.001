.title KiCad schematic
.include "models/AL8805.spice.txt"
.include "models/B260A.spice.txt"
.include "models/C2012X5R1H475K125AB_p.mod"
.include "models/C2012X7R2A104K125AE_p.mod"
.include "models/C2012X7R2E103K125AA_p.mod"
.include "models/C3225X7T2J104M160AC_p.mod"
.include "models/XPE_SPICE.lib"
XU103 /SW 0 /CTRL /A VCC AL8805
XU104 /CTRL 0 C2012X7R2E103K125AA_p
R103 /CTRL /DIMM 1k
XU102 VCC 0 C2012X7R2A104K125AE_p
XU101 VCC 0 C2012X5R1H475K125AB_p
XU105 /A /K C3225X7T2J104M160AC_p
L101 /SW /K 68u rser=0.089
R101 VCC /A {Rs1}
D101 /SW VCC DI_B260A
V101 VCC 0 {VCC}
V102 /DIMM 0 {VDIMM}
R102 VCC /A {Rs2}
D201 /A /LOAD/1 XLampXPEwhite
D202 /LOAD/1 /LOAD/2 XLampXPEwhite
D203 /LOAD/2 /LOAD/3 XLampXPEwhite
D204 /LOAD/3 /LOAD/4 XLampXPEwhite
D205 /LOAD/4 /LOAD/5 XLampXPEwhite
D206 /LOAD/5 /LOAD/6 XLampXPEwhite
D208 /LOAD/7 /K XLampXPEwhite
D207 /LOAD/6 /LOAD/7 XLampXPEwhite
D209 /A /LOAD/1 XLampXPEwhite
D210 /LOAD/1 /LOAD/2 XLampXPEwhite
D211 /LOAD/2 /LOAD/3 XLampXPEwhite
D212 /LOAD/3 /LOAD/4 XLampXPEwhite
D213 /LOAD/4 /LOAD/5 XLampXPEwhite
D214 /LOAD/5 /LOAD/6 XLampXPEwhite
D216 /LOAD/7 /K XLampXPEwhite
D215 /LOAD/6 /LOAD/7 XLampXPEwhite
.end
